`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:07:18 02/26/2014 
// Design Name: 
// Module Name:    arya 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module arya(
    input clk,
    input reset,
    input [9:0] mem_addr_in,
    input [63:0] mem_data_in,
    input debug_on,
    output [63:0] mem_data_out,
    output [9:0] mem_addr_out
    );


endmodule
